`timescale 1ns/1ps
/*
Module Name: 
Language: System Verilog
Author: Justin Killam
Description:

Parameters:


Inputs:


Outputs:


Module Instantiation Skeleton:

*/

module MIPS_Control_Unit (
    input [5:0]opcode,
    input [5:0]funct,
    output RFWE,
    output RFDSel,
    output ALUInSel,
    output Branch,
    output DMWE,
    output MtoRFSel,
    output Jump,
    output [3:0]ALUsel
    );

endmodule